module vffmpeg

// info Prints information
fn info() {
	println('Read the docs, if there ever is any..')
}
