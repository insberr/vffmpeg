module vffmpeg

pub fn (video Video) details() {
	println('video details')
}