module vffmpeg

pub fn split() {
	println('split stuff')
}